(VARIABLE)
d_Linc_to_PAC,int,0x806D1C,
d_CarNum,HEX,0x806D18,
ddddd,int,0x806D1B,
d_CI_Index,int,0x806D17,
d_CI_Fault,int,0x806D16,
d_CarConfig_St,int,0x806D1A,
d_CarConfig,int,0x806D19,
d_MDS_info,HEX,0x806912,
d_MDS_TX_Cnt_A,int,0x806F13,
d_MDS_TX_Cnt_B,int,0x806F14,
m_nDebugCnt,int,0x8071E6,
(ADDRESS)
0x000000,0x0003083A,HEX
(SEPARE ADDRESS)
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
,,
